// problema1.v

// Generated using ACDS version 13.1 162 at 2019.09.14.02:03:27

`timescale 1 ps / 1 ps
module problema1 (
		input  wire       clk_clk,         //      clk.clk
		input  wire       reset_reset_n,   //    reset.reset_n
		output wire [7:0] data_export,     //     data.export
		output wire       enable_export,   //   enable.export
		output wire       rs_export,       //       rs.export
		output wire       rw_export,       //       rw.export
		output wire [9:0] y1_export,       //       y1.export
		output wire [9:0] y2_export,       //       y2.export
		output wire [9:0] xbola_export,    //    xbola.export
		output wire [9:0] ybola_export,    //    ybola.export
		input  wire       endframe_export, // endframe.export
		input  wire [7:0] ad0_export,      //      ad0.export
		input  wire [7:0] ad1_export,      //      ad1.export
		input  wire       adc_busy_export, // adc_busy.export
		input  wire [1:0] button_export    //   button.export
	);

	wire  [31:0] processor_custom_instruction_master_result;                                   // processor_custom_instruction_master_translator:ci_slave_result -> processor:E_ci_result
	wire   [4:0] processor_custom_instruction_master_b;                                        // processor:D_ci_b -> processor_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] processor_custom_instruction_master_c;                                        // processor:D_ci_c -> processor_custom_instruction_master_translator:ci_slave_c
	wire         processor_custom_instruction_master_done;                                     // processor_custom_instruction_master_translator:ci_slave_multi_done -> processor:E_ci_multi_done
	wire         processor_custom_instruction_master_clk_en;                                   // processor:E_ci_multi_clk_en -> processor_custom_instruction_master_translator:ci_slave_multi_clken
	wire   [4:0] processor_custom_instruction_master_a;                                        // processor:D_ci_a -> processor_custom_instruction_master_translator:ci_slave_a
	wire   [7:0] processor_custom_instruction_master_n;                                        // processor:D_ci_n -> processor_custom_instruction_master_translator:ci_slave_n
	wire         processor_custom_instruction_master_writerc;                                  // processor:D_ci_writerc -> processor_custom_instruction_master_translator:ci_slave_writerc
	wire         processor_custom_instruction_master_clk;                                      // processor:E_ci_multi_clock -> processor_custom_instruction_master_translator:ci_slave_multi_clk
	wire         processor_custom_instruction_master_reset_req;                                // processor:E_ci_multi_reset_req -> processor_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         processor_custom_instruction_master_start;                                    // processor:E_ci_multi_start -> processor_custom_instruction_master_translator:ci_slave_multi_start
	wire  [31:0] processor_custom_instruction_master_dataa;                                    // processor:E_ci_dataa -> processor_custom_instruction_master_translator:ci_slave_dataa
	wire         processor_custom_instruction_master_readra;                                   // processor:D_ci_readra -> processor_custom_instruction_master_translator:ci_slave_readra
	wire         processor_custom_instruction_master_reset;                                    // processor:E_ci_multi_reset -> processor_custom_instruction_master_translator:ci_slave_multi_reset
	wire  [31:0] processor_custom_instruction_master_datab;                                    // processor:E_ci_datab -> processor_custom_instruction_master_translator:ci_slave_datab
	wire         processor_custom_instruction_master_readrb;                                   // processor:D_ci_readrb -> processor_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] processor_custom_instruction_master_translator_multi_ci_master_result;        // processor_custom_instruction_master_multi_xconnect:ci_slave_result -> processor_custom_instruction_master_translator:multi_ci_master_result
	wire   [4:0] processor_custom_instruction_master_translator_multi_ci_master_b;             // processor_custom_instruction_master_translator:multi_ci_master_b -> processor_custom_instruction_master_multi_xconnect:ci_slave_b
	wire   [4:0] processor_custom_instruction_master_translator_multi_ci_master_c;             // processor_custom_instruction_master_translator:multi_ci_master_c -> processor_custom_instruction_master_multi_xconnect:ci_slave_c
	wire   [4:0] processor_custom_instruction_master_translator_multi_ci_master_a;             // processor_custom_instruction_master_translator:multi_ci_master_a -> processor_custom_instruction_master_multi_xconnect:ci_slave_a
	wire         processor_custom_instruction_master_translator_multi_ci_master_clk_en;        // processor_custom_instruction_master_translator:multi_ci_master_clken -> processor_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire         processor_custom_instruction_master_translator_multi_ci_master_done;          // processor_custom_instruction_master_multi_xconnect:ci_slave_done -> processor_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] processor_custom_instruction_master_translator_multi_ci_master_n;             // processor_custom_instruction_master_translator:multi_ci_master_n -> processor_custom_instruction_master_multi_xconnect:ci_slave_n
	wire         processor_custom_instruction_master_translator_multi_ci_master_writerc;       // processor_custom_instruction_master_translator:multi_ci_master_writerc -> processor_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         processor_custom_instruction_master_translator_multi_ci_master_clk;           // processor_custom_instruction_master_translator:multi_ci_master_clk -> processor_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         processor_custom_instruction_master_translator_multi_ci_master_reset_req;     // processor_custom_instruction_master_translator:multi_ci_master_reset_req -> processor_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         processor_custom_instruction_master_translator_multi_ci_master_start;         // processor_custom_instruction_master_translator:multi_ci_master_start -> processor_custom_instruction_master_multi_xconnect:ci_slave_start
	wire  [31:0] processor_custom_instruction_master_translator_multi_ci_master_dataa;         // processor_custom_instruction_master_translator:multi_ci_master_dataa -> processor_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         processor_custom_instruction_master_translator_multi_ci_master_readra;        // processor_custom_instruction_master_translator:multi_ci_master_readra -> processor_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire         processor_custom_instruction_master_translator_multi_ci_master_reset;         // processor_custom_instruction_master_translator:multi_ci_master_reset -> processor_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire  [31:0] processor_custom_instruction_master_translator_multi_ci_master_datab;         // processor_custom_instruction_master_translator:multi_ci_master_datab -> processor_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire         processor_custom_instruction_master_translator_multi_ci_master_readrb;        // processor_custom_instruction_master_translator:multi_ci_master_readrb -> processor_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master0_result;         // processor_custom_instruction_master_multi_slave_translator0:ci_slave_result -> processor_custom_instruction_master_multi_xconnect:ci_master0_result
	wire   [4:0] processor_custom_instruction_master_multi_xconnect_ci_master0_b;              // processor_custom_instruction_master_multi_xconnect:ci_master0_b -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire   [4:0] processor_custom_instruction_master_multi_xconnect_ci_master0_c;              // processor_custom_instruction_master_multi_xconnect:ci_master0_c -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_done;           // processor_custom_instruction_master_multi_slave_translator0:ci_slave_done -> processor_custom_instruction_master_multi_xconnect:ci_master0_done
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // processor_custom_instruction_master_multi_xconnect:ci_master0_clken -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [4:0] processor_custom_instruction_master_multi_xconnect_ci_master0_a;              // processor_custom_instruction_master_multi_xconnect:ci_master0_a -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [7:0] processor_custom_instruction_master_multi_xconnect_ci_master0_n;              // processor_custom_instruction_master_multi_xconnect:ci_master0_n -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // processor_custom_instruction_master_multi_xconnect:ci_master0_writerc -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // processor_custom_instruction_master_multi_xconnect:ci_master0_ipending -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_clk;            // processor_custom_instruction_master_multi_xconnect:ci_master0_clk -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // processor_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_start;          // processor_custom_instruction_master_multi_xconnect:ci_master0_start -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // processor_custom_instruction_master_multi_xconnect:ci_master0_dataa -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_readra;         // processor_custom_instruction_master_multi_xconnect:ci_master0_readra -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_reset;          // processor_custom_instruction_master_multi_xconnect:ci_master0_reset -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master0_datab;          // processor_custom_instruction_master_multi_xconnect:ci_master0_datab -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // processor_custom_instruction_master_multi_xconnect:ci_master0_readrb -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire         processor_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // processor_custom_instruction_master_multi_xconnect:ci_master0_estatus -> processor_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire  [31:0] processor_custom_instruction_master_multi_slave_translator0_ci_master_result; // display_0:result -> processor_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         processor_custom_instruction_master_multi_slave_translator0_ci_master_start;  // processor_custom_instruction_master_multi_slave_translator0:ci_master_start -> display_0:iniciar
	wire  [31:0] processor_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // processor_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> display_0:dataA
	wire         processor_custom_instruction_master_multi_slave_translator0_ci_master_done;   // display_0:done -> processor_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         processor_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // processor_custom_instruction_master_multi_slave_translator0:ci_master_clken -> display_0:clk_en
	wire         processor_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // processor_custom_instruction_master_multi_slave_translator0:ci_master_reset -> display_0:reset
	wire  [31:0] processor_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // processor_custom_instruction_master_multi_slave_translator0:ci_master_datab -> display_0:dataB
	wire         processor_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // processor_custom_instruction_master_multi_slave_translator0:ci_master_clk -> display_0:clk
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master1_result;         // processor_custom_instruction_master_multi_slave_translator1:ci_slave_result -> processor_custom_instruction_master_multi_xconnect:ci_master1_result
	wire   [4:0] processor_custom_instruction_master_multi_xconnect_ci_master1_b;              // processor_custom_instruction_master_multi_xconnect:ci_master1_b -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_b
	wire   [4:0] processor_custom_instruction_master_multi_xconnect_ci_master1_c;              // processor_custom_instruction_master_multi_xconnect:ci_master1_c -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_c
	wire         processor_custom_instruction_master_multi_xconnect_ci_master1_done;           // processor_custom_instruction_master_multi_slave_translator1:ci_slave_done -> processor_custom_instruction_master_multi_xconnect:ci_master1_done
	wire         processor_custom_instruction_master_multi_xconnect_ci_master1_clk_en;         // processor_custom_instruction_master_multi_xconnect:ci_master1_clken -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_clken
	wire   [4:0] processor_custom_instruction_master_multi_xconnect_ci_master1_a;              // processor_custom_instruction_master_multi_xconnect:ci_master1_a -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_a
	wire   [7:0] processor_custom_instruction_master_multi_xconnect_ci_master1_n;              // processor_custom_instruction_master_multi_xconnect:ci_master1_n -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_n
	wire         processor_custom_instruction_master_multi_xconnect_ci_master1_writerc;        // processor_custom_instruction_master_multi_xconnect:ci_master1_writerc -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_writerc
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master1_ipending;       // processor_custom_instruction_master_multi_xconnect:ci_master1_ipending -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_ipending
	wire         processor_custom_instruction_master_multi_xconnect_ci_master1_clk;            // processor_custom_instruction_master_multi_xconnect:ci_master1_clk -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_clk
	wire         processor_custom_instruction_master_multi_xconnect_ci_master1_reset_req;      // processor_custom_instruction_master_multi_xconnect:ci_master1_reset_req -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_reset_req
	wire         processor_custom_instruction_master_multi_xconnect_ci_master1_start;          // processor_custom_instruction_master_multi_xconnect:ci_master1_start -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_start
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master1_dataa;          // processor_custom_instruction_master_multi_xconnect:ci_master1_dataa -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_dataa
	wire         processor_custom_instruction_master_multi_xconnect_ci_master1_readra;         // processor_custom_instruction_master_multi_xconnect:ci_master1_readra -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_readra
	wire         processor_custom_instruction_master_multi_xconnect_ci_master1_reset;          // processor_custom_instruction_master_multi_xconnect:ci_master1_reset -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_reset
	wire  [31:0] processor_custom_instruction_master_multi_xconnect_ci_master1_datab;          // processor_custom_instruction_master_multi_xconnect:ci_master1_datab -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_datab
	wire         processor_custom_instruction_master_multi_xconnect_ci_master1_readrb;         // processor_custom_instruction_master_multi_xconnect:ci_master1_readrb -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_readrb
	wire         processor_custom_instruction_master_multi_xconnect_ci_master1_estatus;        // processor_custom_instruction_master_multi_xconnect:ci_master1_estatus -> processor_custom_instruction_master_multi_slave_translator1:ci_slave_estatus
	wire  [31:0] processor_custom_instruction_master_multi_slave_translator1_ci_master_result; // random:result -> processor_custom_instruction_master_multi_slave_translator1:ci_master_result
	wire         processor_custom_instruction_master_multi_slave_translator1_ci_master_start;  // processor_custom_instruction_master_multi_slave_translator1:ci_master_start -> random:start
	wire  [31:0] processor_custom_instruction_master_multi_slave_translator1_ci_master_dataa;  // processor_custom_instruction_master_multi_slave_translator1:ci_master_dataa -> random:dataA
	wire         processor_custom_instruction_master_multi_slave_translator1_ci_master_done;   // random:done -> processor_custom_instruction_master_multi_slave_translator1:ci_master_done
	wire         processor_custom_instruction_master_multi_slave_translator1_ci_master_clk_en; // processor_custom_instruction_master_multi_slave_translator1:ci_master_clken -> random:clk_en
	wire         processor_custom_instruction_master_multi_slave_translator1_ci_master_reset;  // processor_custom_instruction_master_multi_slave_translator1:ci_master_reset -> random:reset
	wire  [31:0] processor_custom_instruction_master_multi_slave_translator1_ci_master_datab;  // processor_custom_instruction_master_multi_slave_translator1:ci_master_datab -> random:dataB
	wire         processor_custom_instruction_master_multi_slave_translator1_ci_master_clk;    // processor_custom_instruction_master_multi_slave_translator1:ci_master_clk -> random:clk
	wire         processor_data_master_waitrequest;                                            // mm_interconnect_0:processor_data_master_waitrequest -> processor:d_waitrequest
	wire  [31:0] processor_data_master_writedata;                                              // processor:d_writedata -> mm_interconnect_0:processor_data_master_writedata
	wire  [13:0] processor_data_master_address;                                                // processor:d_address -> mm_interconnect_0:processor_data_master_address
	wire         processor_data_master_write;                                                  // processor:d_write -> mm_interconnect_0:processor_data_master_write
	wire         processor_data_master_read;                                                   // processor:d_read -> mm_interconnect_0:processor_data_master_read
	wire  [31:0] processor_data_master_readdata;                                               // mm_interconnect_0:processor_data_master_readdata -> processor:d_readdata
	wire         processor_data_master_debugaccess;                                            // processor:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:processor_data_master_debugaccess
	wire   [3:0] processor_data_master_byteenable;                                             // processor:d_byteenable -> mm_interconnect_0:processor_data_master_byteenable
	wire         processor_instruction_master_waitrequest;                                     // mm_interconnect_0:processor_instruction_master_waitrequest -> processor:i_waitrequest
	wire  [13:0] processor_instruction_master_address;                                         // processor:i_address -> mm_interconnect_0:processor_instruction_master_address
	wire         processor_instruction_master_read;                                            // processor:i_read -> mm_interconnect_0:processor_instruction_master_read
	wire  [31:0] processor_instruction_master_readdata;                                        // mm_interconnect_0:processor_instruction_master_readdata -> processor:i_readdata
	wire   [1:0] mm_interconnect_0_button_s1_address;                                          // mm_interconnect_0:button_s1_address -> button:address
	wire  [31:0] mm_interconnect_0_button_s1_readdata;                                         // button:readdata -> mm_interconnect_0:button_s1_readdata
	wire   [1:0] mm_interconnect_0_adc_busy_s1_address;                                        // mm_interconnect_0:ADC_BUSY_s1_address -> ADC_BUSY:address
	wire  [31:0] mm_interconnect_0_adc_busy_s1_readdata;                                       // ADC_BUSY:readdata -> mm_interconnect_0:ADC_BUSY_s1_readdata
	wire  [31:0] mm_interconnect_0_xbola_s1_writedata;                                         // mm_interconnect_0:XBola_s1_writedata -> XBola:writedata
	wire   [1:0] mm_interconnect_0_xbola_s1_address;                                           // mm_interconnect_0:XBola_s1_address -> XBola:address
	wire         mm_interconnect_0_xbola_s1_chipselect;                                        // mm_interconnect_0:XBola_s1_chipselect -> XBola:chipselect
	wire         mm_interconnect_0_xbola_s1_write;                                             // mm_interconnect_0:XBola_s1_write -> XBola:write_n
	wire  [31:0] mm_interconnect_0_xbola_s1_readdata;                                          // XBola:readdata -> mm_interconnect_0:XBola_s1_readdata
	wire   [1:0] mm_interconnect_0_endframe_s1_address;                                        // mm_interconnect_0:endframe_s1_address -> endframe:address
	wire  [31:0] mm_interconnect_0_endframe_s1_readdata;                                       // endframe:readdata -> mm_interconnect_0:endframe_s1_readdata
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                                        // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire   [9:0] mm_interconnect_0_memory_s1_address;                                          // mm_interconnect_0:memory_s1_address -> memory:address
	wire         mm_interconnect_0_memory_s1_chipselect;                                       // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire         mm_interconnect_0_memory_s1_clken;                                            // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire         mm_interconnect_0_memory_s1_write;                                            // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                                         // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                                       // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire  [31:0] mm_interconnect_0_ybola_s1_writedata;                                         // mm_interconnect_0:YBola_s1_writedata -> YBola:writedata
	wire   [1:0] mm_interconnect_0_ybola_s1_address;                                           // mm_interconnect_0:YBola_s1_address -> YBola:address
	wire         mm_interconnect_0_ybola_s1_chipselect;                                        // mm_interconnect_0:YBola_s1_chipselect -> YBola:chipselect
	wire         mm_interconnect_0_ybola_s1_write;                                             // mm_interconnect_0:YBola_s1_write -> YBola:write_n
	wire  [31:0] mm_interconnect_0_ybola_s1_readdata;                                          // YBola:readdata -> mm_interconnect_0:YBola_s1_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                         // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                           // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                             // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                          // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                               // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                                // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                            // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_yplayer1_s1_writedata;                                      // mm_interconnect_0:YPlayer1_s1_writedata -> YPlayer1:writedata
	wire   [1:0] mm_interconnect_0_yplayer1_s1_address;                                        // mm_interconnect_0:YPlayer1_s1_address -> YPlayer1:address
	wire         mm_interconnect_0_yplayer1_s1_chipselect;                                     // mm_interconnect_0:YPlayer1_s1_chipselect -> YPlayer1:chipselect
	wire         mm_interconnect_0_yplayer1_s1_write;                                          // mm_interconnect_0:YPlayer1_s1_write -> YPlayer1:write_n
	wire  [31:0] mm_interconnect_0_yplayer1_s1_readdata;                                       // YPlayer1:readdata -> mm_interconnect_0:YPlayer1_s1_readdata
	wire         mm_interconnect_0_processor_jtag_debug_module_waitrequest;                    // processor:jtag_debug_module_waitrequest -> mm_interconnect_0:processor_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_processor_jtag_debug_module_writedata;                      // mm_interconnect_0:processor_jtag_debug_module_writedata -> processor:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_processor_jtag_debug_module_address;                        // mm_interconnect_0:processor_jtag_debug_module_address -> processor:jtag_debug_module_address
	wire         mm_interconnect_0_processor_jtag_debug_module_write;                          // mm_interconnect_0:processor_jtag_debug_module_write -> processor:jtag_debug_module_write
	wire         mm_interconnect_0_processor_jtag_debug_module_read;                           // mm_interconnect_0:processor_jtag_debug_module_read -> processor:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_processor_jtag_debug_module_readdata;                       // processor:jtag_debug_module_readdata -> mm_interconnect_0:processor_jtag_debug_module_readdata
	wire         mm_interconnect_0_processor_jtag_debug_module_debugaccess;                    // mm_interconnect_0:processor_jtag_debug_module_debugaccess -> processor:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_processor_jtag_debug_module_byteenable;                     // mm_interconnect_0:processor_jtag_debug_module_byteenable -> processor:jtag_debug_module_byteenable
	wire   [1:0] mm_interconnect_0_ad0_s1_address;                                             // mm_interconnect_0:AD0_s1_address -> AD0:address
	wire  [31:0] mm_interconnect_0_ad0_s1_readdata;                                            // AD0:readdata -> mm_interconnect_0:AD0_s1_readdata
	wire   [1:0] mm_interconnect_0_ad1_s1_address;                                             // mm_interconnect_0:AD1_s1_address -> AD1:address
	wire  [31:0] mm_interconnect_0_ad1_s1_readdata;                                            // AD1:readdata -> mm_interconnect_0:AD1_s1_readdata
	wire  [31:0] mm_interconnect_0_yplayer2_s1_writedata;                                      // mm_interconnect_0:YPlayer2_s1_writedata -> YPlayer2:writedata
	wire   [1:0] mm_interconnect_0_yplayer2_s1_address;                                        // mm_interconnect_0:YPlayer2_s1_address -> YPlayer2:address
	wire         mm_interconnect_0_yplayer2_s1_chipselect;                                     // mm_interconnect_0:YPlayer2_s1_chipselect -> YPlayer2:chipselect
	wire         mm_interconnect_0_yplayer2_s1_write;                                          // mm_interconnect_0:YPlayer2_s1_write -> YPlayer2:write_n
	wire  [31:0] mm_interconnect_0_yplayer2_s1_readdata;                                       // YPlayer2:readdata -> mm_interconnect_0:YPlayer2_s1_readdata
	wire         irq_mapper_receiver0_irq;                                                     // jtag:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] processor_d_irq_irq;                                                          // irq_mapper:sender_irq -> processor:d_irq
	wire         rst_controller_reset_out_reset;                                               // rst_controller:reset_out -> [AD0:reset_n, AD1:reset_n, ADC_BUSY:reset_n, XBola:reset_n, YBola:reset_n, YPlayer1:reset_n, YPlayer2:reset_n, button:reset_n, endframe:reset_n, irq_mapper:reset, jtag:rst_n, memory:reset, mm_interconnect_0:processor_reset_n_reset_bridge_in_reset_reset, processor:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                           // rst_controller:reset_req -> [memory:reset_req, processor:reset_req, rst_translator:reset_req_in]
	wire         processor_jtag_debug_module_reset_reset;                                      // processor:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	problema1_processor processor (
		.clk                                   (clk_clk),                                                   //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                           //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                        //                          .reset_req
		.d_address                             (processor_data_master_address),                             //               data_master.address
		.d_byteenable                          (processor_data_master_byteenable),                          //                          .byteenable
		.d_read                                (processor_data_master_read),                                //                          .read
		.d_readdata                            (processor_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (processor_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (processor_data_master_write),                               //                          .write
		.d_writedata                           (processor_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (processor_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (processor_instruction_master_address),                      //        instruction_master.address
		.i_read                                (processor_instruction_master_read),                         //                          .read
		.i_readdata                            (processor_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (processor_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (processor_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (processor_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_processor_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_processor_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_processor_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_processor_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_processor_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_processor_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_processor_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_processor_jtag_debug_module_writedata),   //                          .writedata
		.E_ci_multi_done                       (processor_custom_instruction_master_done),                  // custom_instruction_master.done
		.E_ci_multi_clk_en                     (processor_custom_instruction_master_clk_en),                //                          .clk_en
		.E_ci_multi_start                      (processor_custom_instruction_master_start),                 //                          .start
		.E_ci_result                           (processor_custom_instruction_master_result),                //                          .result
		.D_ci_a                                (processor_custom_instruction_master_a),                     //                          .a
		.D_ci_b                                (processor_custom_instruction_master_b),                     //                          .b
		.D_ci_c                                (processor_custom_instruction_master_c),                     //                          .c
		.D_ci_n                                (processor_custom_instruction_master_n),                     //                          .n
		.D_ci_readra                           (processor_custom_instruction_master_readra),                //                          .readra
		.D_ci_readrb                           (processor_custom_instruction_master_readrb),                //                          .readrb
		.D_ci_writerc                          (processor_custom_instruction_master_writerc),               //                          .writerc
		.E_ci_dataa                            (processor_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_datab                            (processor_custom_instruction_master_datab),                 //                          .datab
		.E_ci_multi_clock                      (processor_custom_instruction_master_clk),                   //                          .clk
		.E_ci_multi_reset                      (processor_custom_instruction_master_reset),                 //                          .reset
		.E_ci_multi_reset_req                  (processor_custom_instruction_master_reset_req)              //                          .reset_req
	);

	problema1_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)      //       .reset_req
	);

	problema1_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	display display_0 (
		.clk     (processor_custom_instruction_master_multi_slave_translator0_ci_master_clk),    // nios_custom_instruction_slave.clk
		.clk_en  (processor_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //                              .clk_en
		.dataA   (processor_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //                              .dataa
		.dataB   (processor_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //                              .datab
		.done    (processor_custom_instruction_master_multi_slave_translator0_ci_master_done),   //                              .done
		.iniciar (processor_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                              .start
		.reset   (processor_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //                              .reset
		.result  (processor_custom_instruction_master_multi_slave_translator0_ci_master_result), //                              .result
		.data    (data_export),                                                                  //                 conduit_end_1.export
		.enable  (enable_export),                                                                //                 conduit_end_2.export
		.rs      (rs_export),                                                                    //                 conduit_end_3.export
		.rw      (rw_export)                                                                     //                 conduit_end_4.export
	);

	problema1_YPlayer1 yplayer1 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_yplayer1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yplayer1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yplayer1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yplayer1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yplayer1_s1_readdata),   //                    .readdata
		.out_port   (y1_export)                                 // external_connection.export
	);

	problema1_YPlayer1 yplayer2 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_yplayer2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yplayer2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yplayer2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yplayer2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yplayer2_s1_readdata),   //                    .readdata
		.out_port   (y2_export)                                 // external_connection.export
	);

	problema1_YPlayer1 xbola (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_xbola_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_xbola_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_xbola_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_xbola_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_xbola_s1_readdata),   //                    .readdata
		.out_port   (xbola_export)                           // external_connection.export
	);

	problema1_YPlayer1 ybola (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_ybola_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ybola_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ybola_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ybola_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ybola_s1_readdata),   //                    .readdata
		.out_port   (ybola_export)                           // external_connection.export
	);

	problema1_endframe endframe (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_endframe_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_endframe_s1_readdata), //                    .readdata
		.in_port  (endframe_export)                         // external_connection.export
	);

	problema1_AD0 ad0 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_ad0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ad0_s1_readdata), //                    .readdata
		.in_port  (ad0_export)                         // external_connection.export
	);

	problema1_AD0 ad1 (
		.clk      (clk_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_ad1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ad1_s1_readdata), //                    .readdata
		.in_port  (ad1_export)                         // external_connection.export
	);

	problema1_endframe adc_busy (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_adc_busy_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_adc_busy_s1_readdata), //                    .readdata
		.in_port  (adc_busy_export)                         // external_connection.export
	);

	random random (
		.clk    (processor_custom_instruction_master_multi_slave_translator1_ci_master_clk),    // nios_custom_instruction_slave.clk
		.clk_en (processor_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //                              .clk_en
		.reset  (processor_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //                              .reset
		.start  (processor_custom_instruction_master_multi_slave_translator1_ci_master_start),  //                              .start
		.dataA  (processor_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  //                              .dataa
		.dataB  (processor_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //                              .datab
		.done   (processor_custom_instruction_master_multi_slave_translator1_ci_master_done),   //                              .done
		.result (processor_custom_instruction_master_multi_slave_translator1_ci_master_result)  //                              .result
	);

	problema1_button button (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_button_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_s1_readdata), //                    .readdata
		.in_port  (button_export)                         // external_connection.export
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) processor_custom_instruction_master_translator (
		.ci_slave_dataa            (processor_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (processor_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (processor_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (processor_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (processor_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (processor_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (processor_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (processor_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (processor_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (processor_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (),                                                                         //                .ipending
		.ci_slave_estatus          (),                                                                         //                .estatus
		.ci_slave_multi_clk        (processor_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (processor_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (processor_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (processor_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (processor_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (processor_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (),                                                                         //  comb_ci_master.dataa
		.comb_ci_master_datab      (),                                                                         //                .datab
		.comb_ci_master_result     (),                                                                         //                .result
		.comb_ci_master_n          (),                                                                         //                .n
		.comb_ci_master_readra     (),                                                                         //                .readra
		.comb_ci_master_readrb     (),                                                                         //                .readrb
		.comb_ci_master_writerc    (),                                                                         //                .writerc
		.comb_ci_master_a          (),                                                                         //                .a
		.comb_ci_master_b          (),                                                                         //                .b
		.comb_ci_master_c          (),                                                                         //                .c
		.comb_ci_master_ipending   (),                                                                         //                .ipending
		.comb_ci_master_estatus    (),                                                                         //                .estatus
		.multi_ci_master_clk       (processor_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (processor_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (processor_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (processor_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (processor_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (processor_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (processor_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (processor_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (processor_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (processor_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (processor_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (processor_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (processor_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (processor_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (processor_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (processor_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                     //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                     //     (terminated)
		.ci_slave_multi_result     (),                                                                         //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                              //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                     //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                     //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                     //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                                 //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                                 //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                                  //     (terminated)
	);

	problema1_processor_custom_instruction_master_multi_xconnect processor_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (processor_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (processor_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (processor_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (processor_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (processor_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (processor_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (processor_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (processor_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (processor_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (processor_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                         //           .ipending
		.ci_slave_estatus     (),                                                                         //           .estatus
		.ci_slave_clk         (processor_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (processor_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (processor_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (processor_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (processor_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (processor_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (processor_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (processor_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (processor_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (processor_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (processor_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (processor_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (processor_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (processor_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (processor_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (processor_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (processor_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (processor_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (processor_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (processor_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (processor_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (processor_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (processor_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (processor_custom_instruction_master_multi_xconnect_ci_master0_done),       //           .done
		.ci_master1_dataa     (processor_custom_instruction_master_multi_xconnect_ci_master1_dataa),      // ci_master1.dataa
		.ci_master1_datab     (processor_custom_instruction_master_multi_xconnect_ci_master1_datab),      //           .datab
		.ci_master1_result    (processor_custom_instruction_master_multi_xconnect_ci_master1_result),     //           .result
		.ci_master1_n         (processor_custom_instruction_master_multi_xconnect_ci_master1_n),          //           .n
		.ci_master1_readra    (processor_custom_instruction_master_multi_xconnect_ci_master1_readra),     //           .readra
		.ci_master1_readrb    (processor_custom_instruction_master_multi_xconnect_ci_master1_readrb),     //           .readrb
		.ci_master1_writerc   (processor_custom_instruction_master_multi_xconnect_ci_master1_writerc),    //           .writerc
		.ci_master1_a         (processor_custom_instruction_master_multi_xconnect_ci_master1_a),          //           .a
		.ci_master1_b         (processor_custom_instruction_master_multi_xconnect_ci_master1_b),          //           .b
		.ci_master1_c         (processor_custom_instruction_master_multi_xconnect_ci_master1_c),          //           .c
		.ci_master1_ipending  (processor_custom_instruction_master_multi_xconnect_ci_master1_ipending),   //           .ipending
		.ci_master1_estatus   (processor_custom_instruction_master_multi_xconnect_ci_master1_estatus),    //           .estatus
		.ci_master1_clk       (processor_custom_instruction_master_multi_xconnect_ci_master1_clk),        //           .clk
		.ci_master1_reset     (processor_custom_instruction_master_multi_xconnect_ci_master1_reset),      //           .reset
		.ci_master1_clken     (processor_custom_instruction_master_multi_xconnect_ci_master1_clk_en),     //           .clk_en
		.ci_master1_reset_req (processor_custom_instruction_master_multi_xconnect_ci_master1_reset_req),  //           .reset_req
		.ci_master1_start     (processor_custom_instruction_master_multi_xconnect_ci_master1_start),      //           .start
		.ci_master1_done      (processor_custom_instruction_master_multi_xconnect_ci_master1_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) processor_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (processor_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (processor_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (processor_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (processor_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (processor_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (processor_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (processor_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (processor_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (processor_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (processor_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (processor_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (processor_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (processor_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (processor_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (processor_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (processor_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (processor_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (processor_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (processor_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (processor_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (processor_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_clk       (processor_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (processor_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (processor_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (processor_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (processor_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_n         (),                                                                             // (terminated)
		.ci_master_readra    (),                                                                             // (terminated)
		.ci_master_readrb    (),                                                                             // (terminated)
		.ci_master_writerc   (),                                                                             // (terminated)
		.ci_master_a         (),                                                                             // (terminated)
		.ci_master_b         (),                                                                             // (terminated)
		.ci_master_c         (),                                                                             // (terminated)
		.ci_master_ipending  (),                                                                             // (terminated)
		.ci_master_estatus   (),                                                                             // (terminated)
		.ci_master_reset_req ()                                                                              // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) processor_custom_instruction_master_multi_slave_translator1 (
		.ci_slave_dataa      (processor_custom_instruction_master_multi_xconnect_ci_master1_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (processor_custom_instruction_master_multi_xconnect_ci_master1_datab),          //          .datab
		.ci_slave_result     (processor_custom_instruction_master_multi_xconnect_ci_master1_result),         //          .result
		.ci_slave_n          (processor_custom_instruction_master_multi_xconnect_ci_master1_n),              //          .n
		.ci_slave_readra     (processor_custom_instruction_master_multi_xconnect_ci_master1_readra),         //          .readra
		.ci_slave_readrb     (processor_custom_instruction_master_multi_xconnect_ci_master1_readrb),         //          .readrb
		.ci_slave_writerc    (processor_custom_instruction_master_multi_xconnect_ci_master1_writerc),        //          .writerc
		.ci_slave_a          (processor_custom_instruction_master_multi_xconnect_ci_master1_a),              //          .a
		.ci_slave_b          (processor_custom_instruction_master_multi_xconnect_ci_master1_b),              //          .b
		.ci_slave_c          (processor_custom_instruction_master_multi_xconnect_ci_master1_c),              //          .c
		.ci_slave_ipending   (processor_custom_instruction_master_multi_xconnect_ci_master1_ipending),       //          .ipending
		.ci_slave_estatus    (processor_custom_instruction_master_multi_xconnect_ci_master1_estatus),        //          .estatus
		.ci_slave_clk        (processor_custom_instruction_master_multi_xconnect_ci_master1_clk),            //          .clk
		.ci_slave_clken      (processor_custom_instruction_master_multi_xconnect_ci_master1_clk_en),         //          .clk_en
		.ci_slave_reset_req  (processor_custom_instruction_master_multi_xconnect_ci_master1_reset_req),      //          .reset_req
		.ci_slave_reset      (processor_custom_instruction_master_multi_xconnect_ci_master1_reset),          //          .reset
		.ci_slave_start      (processor_custom_instruction_master_multi_xconnect_ci_master1_start),          //          .start
		.ci_slave_done       (processor_custom_instruction_master_multi_xconnect_ci_master1_done),           //          .done
		.ci_master_dataa     (processor_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (processor_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //          .datab
		.ci_master_result    (processor_custom_instruction_master_multi_slave_translator1_ci_master_result), //          .result
		.ci_master_clk       (processor_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //          .clk
		.ci_master_clken     (processor_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (processor_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //          .reset
		.ci_master_start     (processor_custom_instruction_master_multi_slave_translator1_ci_master_start),  //          .start
		.ci_master_done      (processor_custom_instruction_master_multi_slave_translator1_ci_master_done),   //          .done
		.ci_master_n         (),                                                                             // (terminated)
		.ci_master_readra    (),                                                                             // (terminated)
		.ci_master_readrb    (),                                                                             // (terminated)
		.ci_master_writerc   (),                                                                             // (terminated)
		.ci_master_a         (),                                                                             // (terminated)
		.ci_master_b         (),                                                                             // (terminated)
		.ci_master_c         (),                                                                             // (terminated)
		.ci_master_ipending  (),                                                                             // (terminated)
		.ci_master_estatus   (),                                                                             // (terminated)
		.ci_master_reset_req ()                                                                              // (terminated)
	);

	problema1_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                 (clk_clk),                                                   //                               clk_0_clk.clk
		.processor_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // processor_reset_n_reset_bridge_in_reset.reset
		.processor_data_master_address                 (processor_data_master_address),                             //                   processor_data_master.address
		.processor_data_master_waitrequest             (processor_data_master_waitrequest),                         //                                        .waitrequest
		.processor_data_master_byteenable              (processor_data_master_byteenable),                          //                                        .byteenable
		.processor_data_master_read                    (processor_data_master_read),                                //                                        .read
		.processor_data_master_readdata                (processor_data_master_readdata),                            //                                        .readdata
		.processor_data_master_write                   (processor_data_master_write),                               //                                        .write
		.processor_data_master_writedata               (processor_data_master_writedata),                           //                                        .writedata
		.processor_data_master_debugaccess             (processor_data_master_debugaccess),                         //                                        .debugaccess
		.processor_instruction_master_address          (processor_instruction_master_address),                      //            processor_instruction_master.address
		.processor_instruction_master_waitrequest      (processor_instruction_master_waitrequest),                  //                                        .waitrequest
		.processor_instruction_master_read             (processor_instruction_master_read),                         //                                        .read
		.processor_instruction_master_readdata         (processor_instruction_master_readdata),                     //                                        .readdata
		.AD0_s1_address                                (mm_interconnect_0_ad0_s1_address),                          //                                  AD0_s1.address
		.AD0_s1_readdata                               (mm_interconnect_0_ad0_s1_readdata),                         //                                        .readdata
		.AD1_s1_address                                (mm_interconnect_0_ad1_s1_address),                          //                                  AD1_s1.address
		.AD1_s1_readdata                               (mm_interconnect_0_ad1_s1_readdata),                         //                                        .readdata
		.ADC_BUSY_s1_address                           (mm_interconnect_0_adc_busy_s1_address),                     //                             ADC_BUSY_s1.address
		.ADC_BUSY_s1_readdata                          (mm_interconnect_0_adc_busy_s1_readdata),                    //                                        .readdata
		.button_s1_address                             (mm_interconnect_0_button_s1_address),                       //                               button_s1.address
		.button_s1_readdata                            (mm_interconnect_0_button_s1_readdata),                      //                                        .readdata
		.endframe_s1_address                           (mm_interconnect_0_endframe_s1_address),                     //                             endframe_s1.address
		.endframe_s1_readdata                          (mm_interconnect_0_endframe_s1_readdata),                    //                                        .readdata
		.jtag_avalon_jtag_slave_address                (mm_interconnect_0_jtag_avalon_jtag_slave_address),          //                  jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_avalon_jtag_slave_write),            //                                        .write
		.jtag_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_avalon_jtag_slave_read),             //                                        .read
		.jtag_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),         //                                        .readdata
		.jtag_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),        //                                        .writedata
		.jtag_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),      //                                        .waitrequest
		.jtag_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),       //                                        .chipselect
		.memory_s1_address                             (mm_interconnect_0_memory_s1_address),                       //                               memory_s1.address
		.memory_s1_write                               (mm_interconnect_0_memory_s1_write),                         //                                        .write
		.memory_s1_readdata                            (mm_interconnect_0_memory_s1_readdata),                      //                                        .readdata
		.memory_s1_writedata                           (mm_interconnect_0_memory_s1_writedata),                     //                                        .writedata
		.memory_s1_byteenable                          (mm_interconnect_0_memory_s1_byteenable),                    //                                        .byteenable
		.memory_s1_chipselect                          (mm_interconnect_0_memory_s1_chipselect),                    //                                        .chipselect
		.memory_s1_clken                               (mm_interconnect_0_memory_s1_clken),                         //                                        .clken
		.processor_jtag_debug_module_address           (mm_interconnect_0_processor_jtag_debug_module_address),     //             processor_jtag_debug_module.address
		.processor_jtag_debug_module_write             (mm_interconnect_0_processor_jtag_debug_module_write),       //                                        .write
		.processor_jtag_debug_module_read              (mm_interconnect_0_processor_jtag_debug_module_read),        //                                        .read
		.processor_jtag_debug_module_readdata          (mm_interconnect_0_processor_jtag_debug_module_readdata),    //                                        .readdata
		.processor_jtag_debug_module_writedata         (mm_interconnect_0_processor_jtag_debug_module_writedata),   //                                        .writedata
		.processor_jtag_debug_module_byteenable        (mm_interconnect_0_processor_jtag_debug_module_byteenable),  //                                        .byteenable
		.processor_jtag_debug_module_waitrequest       (mm_interconnect_0_processor_jtag_debug_module_waitrequest), //                                        .waitrequest
		.processor_jtag_debug_module_debugaccess       (mm_interconnect_0_processor_jtag_debug_module_debugaccess), //                                        .debugaccess
		.XBola_s1_address                              (mm_interconnect_0_xbola_s1_address),                        //                                XBola_s1.address
		.XBola_s1_write                                (mm_interconnect_0_xbola_s1_write),                          //                                        .write
		.XBola_s1_readdata                             (mm_interconnect_0_xbola_s1_readdata),                       //                                        .readdata
		.XBola_s1_writedata                            (mm_interconnect_0_xbola_s1_writedata),                      //                                        .writedata
		.XBola_s1_chipselect                           (mm_interconnect_0_xbola_s1_chipselect),                     //                                        .chipselect
		.YBola_s1_address                              (mm_interconnect_0_ybola_s1_address),                        //                                YBola_s1.address
		.YBola_s1_write                                (mm_interconnect_0_ybola_s1_write),                          //                                        .write
		.YBola_s1_readdata                             (mm_interconnect_0_ybola_s1_readdata),                       //                                        .readdata
		.YBola_s1_writedata                            (mm_interconnect_0_ybola_s1_writedata),                      //                                        .writedata
		.YBola_s1_chipselect                           (mm_interconnect_0_ybola_s1_chipselect),                     //                                        .chipselect
		.YPlayer1_s1_address                           (mm_interconnect_0_yplayer1_s1_address),                     //                             YPlayer1_s1.address
		.YPlayer1_s1_write                             (mm_interconnect_0_yplayer1_s1_write),                       //                                        .write
		.YPlayer1_s1_readdata                          (mm_interconnect_0_yplayer1_s1_readdata),                    //                                        .readdata
		.YPlayer1_s1_writedata                         (mm_interconnect_0_yplayer1_s1_writedata),                   //                                        .writedata
		.YPlayer1_s1_chipselect                        (mm_interconnect_0_yplayer1_s1_chipselect),                  //                                        .chipselect
		.YPlayer2_s1_address                           (mm_interconnect_0_yplayer2_s1_address),                     //                             YPlayer2_s1.address
		.YPlayer2_s1_write                             (mm_interconnect_0_yplayer2_s1_write),                       //                                        .write
		.YPlayer2_s1_readdata                          (mm_interconnect_0_yplayer2_s1_readdata),                    //                                        .readdata
		.YPlayer2_s1_writedata                         (mm_interconnect_0_yplayer2_s1_writedata),                   //                                        .writedata
		.YPlayer2_s1_chipselect                        (mm_interconnect_0_yplayer2_s1_chipselect)                   //                                        .chipselect
	);

	problema1_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (processor_d_irq_irq)             //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                          // reset_in0.reset
		.reset_in1      (processor_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),          // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),      //          .reset_req
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

endmodule
